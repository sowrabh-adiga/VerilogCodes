module fa4b(a,b,cin,s,cout);
input [3:0]a;
input [3:0]b;
input cin;
output [3:0]s;
output cout;
wire c1,c2,c3;
fa f1 (a[0],b[0],cin,s[0],c1);
fa f2 (a[1],b[1],c1,s[1],c2);
fa f3 (a[2],b[2],c2,s[2],c3);
fa f5 (a[3],b[3],c3,s[3],cout);
endmodule // fa4binput a,[3:0]b,cin,output [3:0]s,coutwire c1,c2,c3;
